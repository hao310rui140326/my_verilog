// sim_define.vh
`define TEST_012
// TODO TEST_005 and TEST_007 Error clean

// Number of ports
parameter PORTS = 4;
// Length field width
parameter LEN_WIDTH = 16;
// Tag field width
parameter TAG_WIDTH = 8;

// 88 -> 856
//"INC","DEC","FIX","RAND"
//"INC","DEC","RAND"
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd88 ,16'd88 ,16'd88 ,16'd88 };
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd112,16'd112,16'd112,16'd112};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd113,16'd113,16'd113,16'd113};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd65,16'd1024,16'd128,16'd48};

`ifdef TEST_001
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd588,16'd588,16'd588,16'd588};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd288,16'd288,16'd288,16'd288};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd88 ,16'd88 ,16'd88 ,16'd88 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN   = {16'd48 ,16'd48 ,16'd48 ,16'd48 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_QUEUE_DEPTH = {16'd1,16'd1,16'd1,16'd20};
parameter [PORTS*TAG_WIDTH-1:0]	DEFAULT_TAG_VALUE   = {8'd4,8'd3,8'd2,8'd1};

parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_TEST_MODE = {4'd2,4'd2,4'd2,4'd2};    //"0=INC","1=DEC","2=FIX","3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_CON_TEST_MODE = {4'd0,4'd0,4'd0,4'd0};    //"0=INC","1=DEC",        "3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MIN       = {  16'd48,  16'd48,  16'd48,  16'd48};
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MAX       = {16'd2048,16'd2048,16'd2048,16'd2048};
`endif

`ifdef TEST_002
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd588,16'd588,16'd588,16'd588};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd288,16'd288,16'd288,16'd288};
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd88 ,16'd88 ,16'd88 ,16'd88 };
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN   = {16'd48 ,16'd48 ,16'd48 ,16'd48 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_QUEUE_DEPTH = {16'd1,16'd1,16'd1,16'd20};
parameter [PORTS*TAG_WIDTH-1:0]	DEFAULT_TAG_VALUE   = {8'd4,8'd3,8'd2,8'd1};

parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_TEST_MODE = {4'd2,4'd2,4'd2,4'd2};    //"0=INC","1=DEC","2=FIX","3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_CON_TEST_MODE = {4'd0,4'd0,4'd0,4'd0};    //"0=INC","1=DEC",        "3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MIN       = {  16'd48,  16'd48,  16'd48,  16'd48};
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MAX       = {16'd2048,16'd2048,16'd2048,16'd2048};
`endif

`ifdef TEST_003
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd588,16'd588,16'd588,16'd588};
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd288,16'd288,16'd288,16'd288};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd88 ,16'd88 ,16'd88 ,16'd88 };
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN   = {16'd48 ,16'd48 ,16'd48 ,16'd48 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_QUEUE_DEPTH = {16'd1,16'd1,16'd1,16'd20};
parameter [PORTS*TAG_WIDTH-1:0]	DEFAULT_TAG_VALUE   = {8'd4,8'd3,8'd2,8'd1};

parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_TEST_MODE = {4'd2,4'd2,4'd2,4'd2};    //"0=INC","1=DEC","2=FIX","3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_CON_TEST_MODE = {4'd0,4'd0,4'd0,4'd0};    //"0=INC","1=DEC",        "3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MIN       = {  16'd48,  16'd48,  16'd48,  16'd48};
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MAX       = {16'd2048,16'd2048,16'd2048,16'd2048};
`endif

`ifdef TEST_004
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd588,16'd588,16'd588,16'd588};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd288,16'd288,16'd288,16'd288};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd88 ,16'd88 ,16'd88 ,16'd88 };
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN   = {16'd48 ,16'd48 ,16'd48 ,16'd48 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_QUEUE_DEPTH = {16'd1,16'd1,16'd1,16'd20};
parameter [PORTS*TAG_WIDTH-1:0]	DEFAULT_TAG_VALUE   = {8'd4,8'd3,8'd2,8'd1};

parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_TEST_MODE = {4'd2,4'd2,4'd2,4'd2};    //"0=INC","1=DEC","2=FIX","3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_CON_TEST_MODE = {4'd0,4'd0,4'd0,4'd0};    //"0=INC","1=DEC",        "3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MIN       = {  16'd48,  16'd48,  16'd48,  16'd48};
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MAX       = {16'd2048,16'd2048,16'd2048,16'd2048};
`endif

`ifdef TEST_005
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd588,16'd588,16'd588,16'd588};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd288,16'd288,16'd288,16'd288};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd88 ,16'd88 ,16'd88 ,16'd88 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN   = {16'd48 ,16'd48 ,16'd48 ,16'd48 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_QUEUE_DEPTH = {16'd1,16'd1,16'd1,16'd200};
parameter [PORTS*TAG_WIDTH-1:0]	DEFAULT_TAG_VALUE   = {8'd4,8'd3,8'd2,8'd1};

parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_TEST_MODE = {4'd2,4'd2,4'd2,4'd0};    //"0=INC","1=DEC","2=FIX","3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_CON_TEST_MODE = {4'd0,4'd0,4'd0,4'd0};    //"0=INC","1=DEC",        "3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MIN       = {16'd48  ,16'd48  ,16'd48  ,16'd60  };
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MAX       = {16'd2048,16'd2048,16'd2048,16'd2048};
`endif

`ifdef TEST_006
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd588,16'd588,16'd588,16'd588};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd288,16'd288,16'd288,16'd288};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd88 ,16'd88 ,16'd88 ,16'd88 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN   = {16'd48 ,16'd48 ,16'd48 ,16'd48 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_QUEUE_DEPTH = {16'd1,16'd1,16'd1,16'd200};
parameter [PORTS*TAG_WIDTH-1:0]	DEFAULT_TAG_VALUE   = {8'd4,8'd3,8'd2,8'd1};

parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_TEST_MODE = {4'd2,4'd2,4'd2,4'd1};    //"0=INC","1=DEC","2=FIX","3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_CON_TEST_MODE = {4'd0,4'd0,4'd0,4'd0};    //"0=INC","1=DEC",        "3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MIN       = {16'd48  ,16'd48  ,16'd48  ,16'd60  };
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MAX       = {16'd1048,16'd1048,16'd1048,16'd888};
`endif

`ifdef TEST_007
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd588,16'd588,16'd588,16'd588};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd288,16'd288,16'd288,16'd288};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd88 ,16'd88 ,16'd88 ,16'd88 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN   = {16'd48 ,16'd48 ,16'd48 ,16'd48 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_QUEUE_DEPTH = {16'd1,16'd1,16'd1,16'd200};
parameter [PORTS*TAG_WIDTH-1:0]	DEFAULT_TAG_VALUE   = {8'd4,8'd3,8'd2,8'd1};

parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_TEST_MODE = {4'd2,4'd2,4'd2,4'd1};    //"0=INC","1=DEC","2=FIX","3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_CON_TEST_MODE = {4'd0,4'd0,4'd0,4'd0};    //"0=INC","1=DEC",        "3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MIN       = {16'd48  ,16'd48  ,16'd48  ,16'd60  };
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MAX       = {16'd256 ,16'd256 ,16'd256 ,16'd256 };
`endif

`ifdef TEST_008
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd588,16'd588,16'd588,16'd588};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd288,16'd288,16'd288,16'd288};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd88 ,16'd88 ,16'd88 ,16'd88 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN   = {16'd48 ,16'd48 ,16'd48 ,16'd48 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_QUEUE_DEPTH = {16'd1,16'd1,16'd1,16'd2000};
parameter [PORTS*TAG_WIDTH-1:0]	DEFAULT_TAG_VALUE   = {8'd4,8'd3,8'd2,8'd1};

parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_TEST_MODE = {4'd2,4'd2,4'd2,4'd1};    //"0=INC","1=DEC","2=FIX","3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_CON_TEST_MODE = {4'd0,4'd0,4'd0,4'd0};    //"0=INC","1=DEC",        "3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MIN       = {16'd48  ,16'd48  ,16'd48  ,16'd60  };
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MAX       = {16'd256 ,16'd256 ,16'd256 ,16'd2000 };
`endif

`ifdef TEST_009
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd588,16'd588,16'd588,16'd588};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd288,16'd288,16'd288,16'd288};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd88 ,16'd88 ,16'd88 ,16'd88 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN   = {16'd48 ,16'd48 ,16'd48 ,16'd48 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_QUEUE_DEPTH = {16'd1,16'd1,16'd1,16'd2000};
parameter [PORTS*TAG_WIDTH-1:0]	DEFAULT_TAG_VALUE   = {8'd4,8'd3,8'd2,8'd1};

parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_TEST_MODE = {4'd2,4'd2,4'd2,4'd0};    //"0=INC","1=DEC","2=FIX","3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_CON_TEST_MODE = {4'd0,4'd0,4'd0,4'd1};    //"0=INC","1=DEC",        "3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MIN       = {16'd48  ,16'd48  ,16'd48  ,16'd48  };
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MAX       = {16'd256 ,16'd256 ,16'd256 ,16'd2000 };
`endif

`ifdef TEST_010
// 四队列：其中三个对列固定发送帧长和数量，一个队列帧长在48到2048随机变化，发送个数为200 + 3
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd588,16'd588,16'd588,16'd588};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd288,16'd288,16'd288,16'd288};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd88 ,16'd88 ,16'd88 ,16'd88 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN   = {16'd48 ,16'd48 ,16'd48 ,16'd48 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_QUEUE_DEPTH = {16'd1,16'd1,16'd1,16'd200};
parameter [PORTS*TAG_WIDTH-1:0]	DEFAULT_TAG_VALUE   = {8'd4,8'd3,8'd2,8'd1};

parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_TEST_MODE = {4'd2,4'd2,4'd2,4'd3};    //"0=INC","1=DEC","2=FIX","3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_CON_TEST_MODE = {4'd0,4'd0,4'd0,4'd3};    //"0=INC","1=DEC",        "3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MIN       = {16'd48  ,16'd48  ,16'd48  ,16'd48  };
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MAX       = {16'd256 ,16'd256 ,16'd256 ,16'd2048};
`endif

`ifdef TEST_011
// 四队列：每队列帧长在48到2048随机变化，发送个数为200*4
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd588,16'd588,16'd588,16'd588};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd288,16'd288,16'd288,16'd288};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd88 ,16'd88 ,16'd88 ,16'd88 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN   = {16'd48 ,16'd48 ,16'd48 ,16'd48 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_QUEUE_DEPTH = {16'd200,16'd200,16'd200,16'd200};
parameter [PORTS*TAG_WIDTH-1:0]	DEFAULT_TAG_VALUE   = {8'd4,8'd3,8'd2,8'd1};

parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_TEST_MODE = {4'd3,4'd3,4'd3,4'd3};    //"0=INC","1=DEC","2=FIX","3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_CON_TEST_MODE = {4'd3,4'd3,4'd3,4'd3};    //"0=INC","1=DEC",        "3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MIN       = {16'd48  ,16'd48  ,16'd48  ,16'd48  };
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MAX       = {16'd256 ,16'd1024,16'd512 ,16'd2048};
`endif

`ifdef TEST_012
// 四队列：每队列帧长在48到1048递增，发送个数为1020*4
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd588,16'd588,16'd588,16'd588};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd288,16'd288,16'd288,16'd288};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd88 ,16'd88 ,16'd88 ,16'd88 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN   = {16'd48 ,16'd48 ,16'd48 ,16'd48 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_QUEUE_DEPTH = {16'd1020,16'd1020,16'd1020,16'd1020};
parameter [PORTS*TAG_WIDTH-1:0]	DEFAULT_TAG_VALUE   = {8'd4,8'd3,8'd2,8'd1};

parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_TEST_MODE = {4'd0,4'd0,4'd0,4'd0};    //"0=INC","1=DEC","2=FIX","3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_CON_TEST_MODE = {4'd3,4'd3,4'd3,4'd3};    //"0=INC","1=DEC",        "3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MIN       = {16'd48  ,16'd48  ,16'd48  ,16'd48  };
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MAX       = {16'd1048 ,16'd1048 ,16'd1048 ,16'd1048};
`endif

`ifdef TEST_013
// 四队列：每队列帧长在1048到2048递增，发送个数为1020*4
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd588,16'd588,16'd588,16'd588};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd288,16'd288,16'd288,16'd288};
//parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN = {16'd88 ,16'd88 ,16'd88 ,16'd88 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_FRAME_LEN   = {16'd48 ,16'd48 ,16'd48 ,16'd48 };
parameter [PORTS*LEN_WIDTH-1:0]	DEFAULT_QUEUE_DEPTH = {16'd1020,16'd1020,16'd1020,16'd1020};
parameter [PORTS*TAG_WIDTH-1:0]	DEFAULT_TAG_VALUE   = {8'd4,8'd3,8'd2,8'd1};

parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_TEST_MODE = {4'd0,4'd0,4'd0,4'd0};    //"0=INC","1=DEC","2=FIX","3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_CON_TEST_MODE = {4'd3,4'd3,4'd3,4'd3};    //"0=INC","1=DEC",        "3=RAND"
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MIN       = {16'd1048 ,16'd1048 ,16'd1048 ,16'd1048};
parameter [PORTS*LEN_WIDTH-1:0] DEFAULT_FRAME_LEN_MAX       = {16'd2048 ,16'd2048 ,16'd2048 ,16'd2048};
`endif
